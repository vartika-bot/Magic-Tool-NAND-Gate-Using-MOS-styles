magic
tech scmos
timestamp 1646421470
<< nwell >>
rect -42 -1 -17 23
rect -7 -3 18 21
rect 68 -4 93 20
rect -9 -39 16 -15
rect 25 -39 50 -15
<< polysilicon >>
rect -31 24 82 27
rect -31 21 -28 24
rect 79 18 82 24
rect -31 -2 -28 1
rect 4 -4 7 -1
rect -8 -11 39 -8
rect 36 -17 39 -11
rect 59 -13 83 -10
rect 80 -16 83 -13
rect 80 -46 83 -34
rect -31 -72 -11 -69
rect 4 -70 7 -67
rect -31 -73 -28 -72
rect -14 -74 -11 -72
rect -14 -77 53 -74
rect 50 -94 53 -77
rect 80 -94 83 -91
rect 50 -97 83 -94
<< ndiffusion >>
rect -39 -17 -20 -14
rect -39 -21 -37 -17
rect -33 -21 -31 -17
rect -39 -24 -31 -21
rect -39 -28 -37 -24
rect -33 -28 -31 -24
rect -39 -30 -31 -28
rect -28 -21 -26 -17
rect -22 -21 -20 -17
rect -28 -24 -20 -21
rect -28 -28 -26 -24
rect -22 -28 -20 -24
rect -28 -30 -20 -28
rect -39 -33 -20 -30
rect 71 -19 80 -16
rect 71 -23 74 -19
rect 78 -23 80 -19
rect 71 -26 80 -23
rect 71 -30 74 -26
rect 78 -30 80 -26
rect 71 -34 80 -30
rect 83 -19 92 -16
rect 83 -23 85 -19
rect 89 -23 92 -19
rect 83 -26 92 -23
rect 83 -30 85 -26
rect 89 -30 92 -26
rect 83 -34 92 -30
rect -39 -43 -20 -40
rect -39 -47 -37 -43
rect -33 -47 -31 -43
rect -39 -50 -31 -47
rect -39 -54 -37 -50
rect -33 -54 -31 -50
rect -39 -56 -31 -54
rect -28 -47 -26 -43
rect -22 -47 -20 -43
rect -28 -50 -20 -47
rect 72 -48 80 -46
rect -28 -54 -26 -50
rect -22 -54 -20 -50
rect -28 -56 -20 -54
rect -39 -59 -20 -56
rect -5 -51 16 -48
rect -5 -55 -2 -51
rect 2 -55 4 -51
rect -5 -59 4 -55
rect -5 -63 -2 -59
rect 2 -63 4 -59
rect -5 -67 4 -63
rect 7 -55 9 -51
rect 13 -55 16 -51
rect 7 -59 16 -55
rect 7 -63 9 -59
rect 13 -63 16 -59
rect 7 -67 16 -63
rect 72 -52 74 -48
rect 78 -52 80 -48
rect 72 -55 80 -52
rect 72 -59 74 -55
rect 78 -59 80 -55
rect 72 -60 80 -59
rect 83 -48 93 -46
rect 83 -52 85 -48
rect 89 -52 93 -48
rect 83 -55 93 -52
rect 83 -59 85 -55
rect 89 -59 93 -55
rect 83 -60 93 -59
rect 72 -64 93 -60
rect -39 -76 -31 -73
rect -39 -80 -37 -76
rect -33 -80 -31 -76
rect -39 -83 -31 -80
rect -39 -87 -37 -83
rect -33 -87 -31 -83
rect -39 -90 -31 -87
rect -28 -76 -20 -73
rect -28 -80 -26 -76
rect -22 -80 -20 -76
rect -28 -83 -20 -80
rect -28 -87 -26 -83
rect -22 -87 -20 -83
rect -28 -90 -20 -87
rect -39 -93 -20 -90
rect 72 -76 93 -73
rect 72 -80 74 -76
rect 78 -80 80 -76
rect 72 -83 80 -80
rect 72 -87 74 -83
rect 78 -87 80 -83
rect 72 -91 80 -87
rect 83 -80 85 -76
rect 89 -80 93 -76
rect 83 -83 93 -80
rect 83 -87 85 -83
rect 89 -87 93 -83
rect 83 -91 93 -87
<< pdiffusion >>
rect -40 18 -31 21
rect -40 14 -37 18
rect -33 14 -31 18
rect -40 9 -31 14
rect -40 5 -37 9
rect -33 5 -31 9
rect -40 1 -31 5
rect -28 18 -19 21
rect -28 14 -26 18
rect -22 14 -19 18
rect -28 9 -19 14
rect -28 5 -26 9
rect -22 5 -19 9
rect -28 1 -19 5
rect -5 16 16 19
rect -5 12 -2 16
rect 2 12 4 16
rect -5 9 4 12
rect -5 5 -2 9
rect 2 5 4 9
rect -5 -1 4 5
rect 7 12 9 16
rect 13 12 16 16
rect 7 9 16 12
rect 7 5 9 9
rect 13 5 16 9
rect 7 -1 16 5
rect 70 16 79 18
rect 70 12 73 16
rect 77 12 79 16
rect 70 9 79 12
rect 70 5 73 9
rect 77 5 79 9
rect 70 3 79 5
rect 82 16 91 18
rect 82 12 84 16
rect 88 12 91 16
rect 82 9 91 12
rect 82 5 84 9
rect 88 5 91 9
rect 82 3 91 5
rect 70 -2 91 3
rect -7 -20 14 -17
rect -7 -24 -4 -20
rect 0 -24 2 -20
rect -7 -27 2 -24
rect -7 -31 -4 -27
rect 0 -31 2 -27
rect -7 -34 2 -31
rect 5 -24 7 -20
rect 11 -24 14 -20
rect 5 -27 14 -24
rect 5 -31 7 -27
rect 11 -31 14 -27
rect 5 -34 14 -31
rect -7 -37 14 -34
rect 27 -20 36 -17
rect 27 -24 30 -20
rect 34 -24 36 -20
rect 27 -27 36 -24
rect 27 -31 30 -27
rect 34 -31 36 -27
rect 27 -34 36 -31
rect 39 -20 48 -17
rect 39 -24 41 -20
rect 45 -24 48 -20
rect 39 -27 48 -24
rect 39 -31 41 -27
rect 45 -31 48 -27
rect 39 -34 48 -31
rect 27 -37 48 -34
<< metal1 >>
rect -37 32 -33 35
rect -37 28 77 32
rect -37 18 -33 28
rect -37 9 -33 14
rect -37 2 -33 5
rect -26 18 -22 19
rect -26 9 -22 14
rect -26 -7 -22 5
rect -2 16 2 28
rect -2 9 2 12
rect -2 1 2 5
rect 9 16 13 18
rect 9 9 13 12
rect -37 -11 -12 -7
rect 9 -9 13 5
rect 73 16 77 28
rect 73 9 77 12
rect 73 2 77 5
rect 84 9 88 12
rect 84 -7 88 5
rect -37 -17 -33 -11
rect -4 -13 34 -9
rect -37 -24 -33 -21
rect -37 -31 -33 -28
rect -26 -17 -22 -16
rect -26 -24 -22 -21
rect -26 -35 -22 -28
rect -4 -20 0 -13
rect -4 -27 0 -24
rect -4 -35 0 -31
rect 7 -20 11 -18
rect 7 -27 11 -24
rect -37 -39 -22 -35
rect -37 -43 -33 -39
rect 7 -43 11 -31
rect 30 -20 34 -13
rect 30 -27 34 -24
rect 30 -35 34 -31
rect 41 -20 45 -18
rect 41 -27 45 -24
rect 41 -43 45 -31
rect 55 -43 59 -13
rect 74 -11 102 -7
rect 74 -19 78 -11
rect 74 -26 78 -23
rect 74 -32 78 -30
rect 85 -19 89 -18
rect 85 -26 89 -23
rect 85 -38 89 -30
rect -37 -50 -33 -47
rect -37 -55 -33 -54
rect -26 -50 -22 -47
rect -26 -64 -22 -54
rect -37 -68 -22 -64
rect -2 -47 59 -43
rect 74 -42 89 -38
rect -2 -51 2 -47
rect 74 -48 78 -42
rect -2 -59 2 -55
rect -2 -65 2 -63
rect 9 -51 13 -50
rect 9 -59 13 -55
rect 74 -55 78 -52
rect 74 -61 78 -59
rect 85 -55 89 -52
rect -37 -76 -33 -68
rect 9 -71 13 -63
rect 85 -66 89 -59
rect 74 -70 89 -66
rect -37 -83 -33 -80
rect -37 -91 -33 -87
rect -26 -76 -22 -75
rect -26 -83 -22 -80
rect -26 -96 -22 -87
rect 74 -76 78 -70
rect 74 -83 78 -80
rect 74 -89 78 -87
rect 85 -76 89 -75
rect 85 -83 89 -80
rect 85 -95 89 -87
<< ntransistor >>
rect -31 -30 -28 -17
rect 80 -34 83 -16
rect -31 -56 -28 -43
rect 4 -67 7 -51
rect 80 -60 83 -46
rect -31 -90 -28 -73
rect 80 -91 83 -76
<< ptransistor >>
rect -31 1 -28 21
rect 4 -1 7 16
rect 79 3 82 18
rect 2 -34 5 -20
rect 36 -34 39 -17
<< polycontact >>
rect -12 -11 -8 -7
rect 55 -13 59 -9
<< ndcontact >>
rect -37 -21 -33 -17
rect -37 -28 -33 -24
rect -26 -21 -22 -17
rect -26 -28 -22 -24
rect 74 -23 78 -19
rect 74 -30 78 -26
rect 85 -23 89 -19
rect 85 -30 89 -26
rect -37 -47 -33 -43
rect -37 -54 -33 -50
rect -26 -47 -22 -43
rect -26 -54 -22 -50
rect -2 -55 2 -51
rect -2 -63 2 -59
rect 9 -55 13 -51
rect 9 -63 13 -59
rect 74 -52 78 -48
rect 74 -59 78 -55
rect 85 -52 89 -48
rect 85 -59 89 -55
rect -37 -80 -33 -76
rect -37 -87 -33 -83
rect -26 -80 -22 -76
rect -26 -87 -22 -83
rect 74 -80 78 -76
rect 74 -87 78 -83
rect 85 -80 89 -76
rect 85 -87 89 -83
<< pdcontact >>
rect -37 14 -33 18
rect -37 5 -33 9
rect -26 14 -22 18
rect -26 5 -22 9
rect -2 12 2 16
rect -2 5 2 9
rect 9 12 13 16
rect 9 5 13 9
rect 73 12 77 16
rect 73 5 77 9
rect 84 12 88 16
rect 84 5 88 9
rect -4 -24 0 -20
rect -4 -31 0 -27
rect 7 -24 11 -20
rect 7 -31 11 -27
rect 30 -24 34 -20
rect 30 -31 34 -27
rect 41 -24 45 -20
rect 41 -31 45 -27
<< labels >>
rlabel metal1 -35 34 -35 34 5 vdd
rlabel polysilicon -30 0 -30 0 1 a
rlabel ntransistor -30 -29 -30 -29 1 c
rlabel ntransistor -30 -55 -30 -55 1 d
rlabel ntransistor -30 -89 -30 -89 1 b
rlabel metal1 -24 -95 -24 -95 1 vss
rlabel polysilicon 5 -2 5 -2 1 ~b
rlabel polysilicon 5 -69 5 -69 1 ~a
rlabel metal1 11 -70 11 -70 1 vss
rlabel metal1 87 -93 87 -93 1 vss
rlabel metal1 100 -9 100 -9 7 output
<< end >>
