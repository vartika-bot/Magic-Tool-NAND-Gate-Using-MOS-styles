magic
tech scmos
timestamp 1646242863
<< nwell >>
rect -35 2 -10 25
rect 2 2 27 25
rect -16 -37 7 -14
<< polysilicon >>
rect 12 27 34 30
rect 12 23 15 27
rect -25 1 -22 4
rect -41 -2 -22 1
rect 12 -2 15 4
rect -35 -71 -32 -2
rect -6 -39 -3 -35
rect -6 -66 -3 -64
rect -35 -74 -3 -71
rect -6 -75 -3 -74
rect -6 -94 -3 -92
rect 29 -100 32 27
rect -6 -102 32 -100
rect 5 -103 32 -102
rect -6 -122 -3 -119
<< ndiffusion >>
rect -14 -50 5 -47
rect -14 -54 -12 -50
rect -8 -54 -6 -50
rect -14 -57 -6 -54
rect -14 -61 -12 -57
rect -8 -61 -6 -57
rect -14 -64 -6 -61
rect -3 -54 -1 -50
rect 3 -54 5 -50
rect -3 -57 5 -54
rect -3 -61 -1 -57
rect 3 -61 5 -57
rect -3 -64 5 -61
rect -14 -78 -6 -75
rect -14 -82 -12 -78
rect -8 -82 -6 -78
rect -14 -85 -6 -82
rect -14 -89 -12 -85
rect -8 -89 -6 -85
rect -14 -92 -6 -89
rect -3 -78 5 -75
rect -3 -82 -1 -78
rect 3 -82 5 -78
rect -3 -85 5 -82
rect -3 -89 -1 -85
rect 3 -89 5 -85
rect -3 -92 5 -89
rect -14 -105 -6 -102
rect -14 -109 -12 -105
rect -8 -109 -6 -105
rect -14 -112 -6 -109
rect -14 -116 -12 -112
rect -8 -116 -6 -112
rect -14 -119 -6 -116
rect -3 -105 5 -103
rect -3 -109 -1 -105
rect 3 -109 5 -105
rect -3 -112 5 -109
rect -3 -116 -1 -112
rect 3 -116 5 -112
rect -3 -119 5 -116
<< pdiffusion >>
rect -33 20 -12 23
rect -33 16 -31 20
rect -27 16 -25 20
rect -33 12 -25 16
rect -33 8 -31 12
rect -27 8 -25 12
rect -33 4 -25 8
rect -22 16 -19 20
rect -15 16 -12 20
rect -22 12 -12 16
rect -22 8 -19 12
rect -15 8 -12 12
rect -22 4 -12 8
rect 4 20 12 23
rect 4 16 6 20
rect 10 16 12 20
rect 4 12 12 16
rect 4 8 6 12
rect 10 8 12 12
rect 4 4 12 8
rect 15 20 25 23
rect 15 16 17 20
rect 21 16 25 20
rect 15 12 25 16
rect 15 8 17 12
rect 21 8 25 12
rect 15 4 25 8
rect -14 -19 5 -16
rect -14 -23 -12 -19
rect -8 -23 -6 -19
rect -14 -26 -6 -23
rect -14 -30 -12 -26
rect -8 -30 -6 -26
rect -14 -35 -6 -30
rect -3 -23 -1 -19
rect 3 -23 5 -19
rect -3 -26 5 -23
rect -3 -30 -1 -26
rect 3 -30 5 -26
rect -3 -35 5 -30
<< metal1 >>
rect -31 31 -27 34
rect -31 27 10 31
rect -31 20 -27 27
rect -31 12 -27 16
rect -31 6 -27 8
rect -19 20 -15 21
rect -19 12 -15 16
rect -19 -4 -15 8
rect 6 20 10 27
rect 6 12 10 16
rect 6 6 10 8
rect 17 20 21 21
rect 17 12 21 16
rect 17 -4 21 8
rect -19 -8 21 -4
rect -12 -19 -8 -8
rect -12 -26 -8 -23
rect -12 -34 -8 -30
rect -1 -19 3 -18
rect -1 -26 3 -23
rect -1 -41 3 -30
rect -12 -45 50 -41
rect -12 -50 -8 -45
rect -12 -57 -8 -54
rect -12 -62 -8 -61
rect -1 -50 3 -49
rect -1 -57 3 -54
rect -1 -68 3 -61
rect -12 -72 3 -68
rect -12 -78 -8 -72
rect -12 -85 -8 -82
rect -12 -90 -8 -89
rect -1 -78 3 -77
rect -1 -85 3 -82
rect -1 -96 3 -89
rect -12 -100 3 -96
rect -12 -105 -8 -100
rect -12 -112 -8 -109
rect -12 -117 -8 -116
rect -1 -105 3 -104
rect -1 -112 3 -109
rect -1 -126 3 -116
<< ntransistor >>
rect -6 -64 -3 -50
rect -6 -92 -3 -75
rect -6 -103 5 -102
rect -6 -119 -3 -103
<< ptransistor >>
rect -25 4 -22 20
rect 12 4 15 23
rect -6 -35 -3 -19
<< ndcontact >>
rect -12 -54 -8 -50
rect -12 -61 -8 -57
rect -1 -54 3 -50
rect -1 -61 3 -57
rect -12 -82 -8 -78
rect -12 -89 -8 -85
rect -1 -82 3 -78
rect -1 -89 3 -85
rect -12 -109 -8 -105
rect -12 -116 -8 -112
rect -1 -109 3 -105
rect -1 -116 3 -112
<< pdcontact >>
rect -31 16 -27 20
rect -31 8 -27 12
rect -19 16 -15 20
rect -19 8 -15 12
rect 6 16 10 20
rect 6 8 10 12
rect 17 16 21 20
rect 17 8 21 12
rect -12 -23 -8 -19
rect -12 -30 -8 -26
rect -1 -23 3 -19
rect -1 -30 3 -26
<< labels >>
rlabel metal1 -29 31 -29 31 5 vdd
rlabel metal1 47 -43 47 -43 7 vdd
<< end >>
