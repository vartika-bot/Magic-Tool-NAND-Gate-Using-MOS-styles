magic
tech scmos
timestamp 1643046998
<< nwell >>
rect -32 -2 -9 12
rect 35 -6 58 9
rect -32 -38 -9 -24
<< polysilicon >>
rect 24 12 75 15
rect -22 -3 -19 1
rect 6 0 9 3
rect 6 -3 21 0
rect -41 -6 -19 -3
rect -22 -12 -19 -6
rect -22 -15 9 -12
rect 6 -23 9 -15
rect 6 -35 9 -32
rect -22 -45 -19 -35
rect 18 -45 21 -3
rect 24 -8 27 12
rect 45 6 48 12
rect 72 8 75 12
rect -40 -48 21 -45
<< ndiffusion >>
rect 0 9 15 12
rect 0 4 1 9
rect 5 4 6 9
rect 0 3 6 4
rect 9 4 10 9
rect 14 4 15 9
rect 9 3 15 4
rect 0 -26 6 -23
rect 0 -31 1 -26
rect 5 -31 6 -26
rect 0 -32 6 -31
rect 9 -26 15 -23
rect 9 -31 10 -26
rect 14 -31 15 -26
rect 9 -32 15 -31
rect 66 7 72 8
rect 66 2 67 7
rect 71 2 72 7
rect 75 7 81 8
rect 75 2 76 7
rect 80 2 81 7
rect 66 -1 81 2
<< pdiffusion >>
rect -29 6 -12 9
rect -29 1 -27 6
rect -23 1 -22 6
rect -19 1 -18 6
rect -14 1 -12 6
rect -29 -30 -12 -27
rect -29 -35 -27 -30
rect -23 -35 -22 -30
rect -19 -35 -18 -30
rect -14 -35 -12 -30
rect 38 5 45 6
rect 38 0 40 5
rect 44 0 45 5
rect 48 5 55 6
rect 48 0 49 5
rect 53 0 55 5
rect 38 -3 55 0
<< metal1 >>
rect -41 16 5 20
rect -41 -6 -37 16
rect -27 6 -23 16
rect 1 9 5 16
rect -18 6 -14 7
rect -18 -5 -14 1
rect 10 -5 14 4
rect 40 5 44 8
rect 76 7 80 13
rect 40 -2 44 0
rect -18 -9 27 -5
rect -40 -20 5 -16
rect -40 -48 -36 -20
rect -27 -30 -23 -20
rect 1 -26 5 -20
rect -18 -30 -14 -29
rect 10 -26 14 -24
rect -18 -40 -14 -35
rect 10 -40 14 -31
rect 23 -40 27 -9
rect 49 -7 53 0
rect 67 -7 71 2
rect 76 0 80 2
rect 49 -11 81 -7
rect -18 -44 27 -40
<< ntransistor >>
rect 6 3 9 9
rect 6 -32 9 -23
rect 72 2 75 8
<< ptransistor >>
rect -22 1 -19 6
rect -22 -35 -19 -30
rect 45 0 48 6
<< ndcontact >>
rect 1 4 5 9
rect 10 4 14 9
rect 1 -31 5 -26
rect 10 -31 14 -26
rect 67 2 71 7
rect 76 2 80 7
<< pdcontact >>
rect -27 1 -23 6
rect -18 1 -14 6
rect -27 -35 -23 -30
rect -18 -35 -14 -30
rect 40 0 44 5
rect 49 0 53 5
<< labels >>
rlabel metal1 79 -9 79 -9 7 out
rlabel polysilicon 46 11 46 11 1 vdd
rlabel metal1 -39 -5 -39 -5 3 a
rlabel metal1 -38 -47 -38 -47 2 b
rlabel metal1 78 10 78 10 7 gnd
<< end >>
