magic
tech scmos
timestamp 1632300303
<< error_p >>
rect -3 12 -2 17
rect -5 10 -2 12
rect -1 11 1 13
rect 2 10 4 12
rect -3 8 -1 10
rect 4 8 6 10
rect -5 7 -2 8
rect 2 7 5 8
rect -3 5 -1 7
rect 4 5 6 7
rect 4 -2 5 5
rect -2 -3 2 -2
rect 4 -3 9 -2
rect -2 -5 -1 -3
rect 1 -7 2 -5
rect 0 -8 8 -7
rect -1 -9 8 -8
rect -1 -10 2 -9
rect 6 -10 9 -9
rect 1 -12 3 -10
rect 8 -12 10 -10
rect -1 -13 2 -12
rect 6 -13 9 -12
rect 1 -15 3 -13
rect 8 -15 10 -13
rect 1 -16 2 -15
rect -2 -22 6 -21
rect 8 -22 9 -15
rect -2 -24 -1 -22
rect 1 -25 2 -24
rect 0 -26 8 -25
rect -1 -27 8 -26
rect -1 -28 2 -27
rect 6 -28 8 -27
rect 1 -30 3 -28
rect 8 -30 10 -28
rect -1 -31 2 -30
rect 6 -31 9 -30
rect 1 -33 3 -31
rect 8 -33 10 -31
<< nwell >>
rect -9 2 8 13
<< polysilicon >>
rect -1 0 1 4
rect -13 -2 1 0
rect 3 -21 5 -16
rect 3 -39 5 -34
<< ndiffusion >>
rect -2 -10 9 -9
rect -2 -12 -1 -10
rect 1 -12 3 -10
rect -2 -13 3 -12
rect -2 -15 -1 -13
rect 1 -15 3 -13
rect -2 -16 3 -15
rect 5 -12 6 -10
rect 8 -12 9 -10
rect 5 -13 9 -12
rect 5 -15 6 -13
rect 8 -15 9 -13
rect 5 -16 9 -15
rect -2 -28 9 -27
rect -2 -30 -1 -28
rect 1 -30 3 -28
rect -2 -31 3 -30
rect -2 -33 -1 -31
rect 1 -33 3 -31
rect -2 -34 3 -33
rect 5 -30 6 -28
rect 8 -30 9 -28
rect 5 -31 9 -30
rect 5 -33 6 -31
rect 8 -33 9 -31
rect 5 -34 9 -33
<< pdiffusion >>
rect -6 10 5 11
rect -6 8 -5 10
rect -3 8 -1 10
rect -6 7 -1 8
rect -6 5 -5 7
rect -3 5 -1 7
rect -6 4 -1 5
rect 1 8 2 10
rect 4 8 5 10
rect 1 7 5 8
rect 1 5 2 7
rect 4 5 5 7
rect 1 4 5 5
<< metal1 >>
rect -5 10 -3 17
rect -5 7 -3 8
rect 2 7 4 8
rect 2 -3 4 5
rect -1 -5 9 -3
rect -1 -10 1 -5
rect -1 -13 1 -12
rect -1 -16 1 -15
rect 6 -10 8 -9
rect 6 -13 8 -12
rect 6 -22 8 -15
rect -1 -24 8 -22
rect -1 -28 1 -24
rect -1 -31 1 -30
rect 6 -31 8 -30
<< ntransistor >>
rect 3 -16 5 -10
rect 3 -34 5 -28
<< ptransistor >>
rect -1 4 1 10
<< ndcontact >>
rect -1 -12 1 -10
rect -1 -15 1 -13
rect 6 -12 8 -10
rect 6 -15 8 -13
rect -1 -30 1 -28
rect -1 -33 1 -31
rect 6 -30 8 -28
rect 6 -33 8 -31
<< pdcontact >>
rect -5 8 -3 10
rect -5 5 -3 7
rect 2 8 4 10
rect 2 5 4 7
<< labels >>
rlabel polysilicon 4 -20 4 -20 1 a
rlabel polysilicon 4 -38 4 -38 1 b
rlabel polysilicon -11 -1 -11 -1 3 gnd
rlabel metal1 -4 16 -4 16 5 vdd
rlabel metal1 6 -4 6 -4 7 out
<< end >>
